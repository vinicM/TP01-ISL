module display (
    input c1,
    input c2,
    input c3,
    input c4,
    input c6,


    output A,
    output B,
    output C,
    output D,
    output E,
    output F,
    output G
);
    
assign A = (((~c1)&(~c2)&(~c3)&(~c4)&(~c6))| ((c1)&(c2)&(c3)&(c4)&(c6)) | ((c2)&(c3)&(~c4)&(~c6)) | ((~c1)&(~c2)&(c4)&(c6)) | ((~c1)&(c3)&(~c4)&(c6)) | ((~c1)&(c3)&(c4)&(~c6)) | ((c1)&(c2)&(~c3)&(~c4)) | ((c1)&(~c2)&(c3)&(~c4)) | ((c1)&(~c2)&(~c3)&(c6)) | ((c1)&(~c2)&(c4)&(~c6)) | ((c2)&(~c3)&(c4)&(~c6)));

assign B = ((c2) | ((~c2)&(c3)) | ((~c2)&(~c3)&(c4)&(c6)) | ((~c2)&(~c3)&(c4)) | ((c1)&(~c2)&(~c3)&(~c4)&(~c6)));

assign C = (((~c2)&(~c4)&(~c6)) | ((~c1)&(~c4)&(~c6)) | ((~c2)&(~c3)&(~c4)&(c6)) | ((~c1)&(~c2)&(~c3)&(c6)) | ((~c1)&(~c2)&(c4)&(~c6)) | ((c1)&(~c2)&(~c3)&(~c4)) | ((c2)&(~c3)&(~c4)&(~c6)) | ((~c1)&(~c2)&(~c4)&(c6)) | ((~c1)&(~c3)&(~c4)&(c6)) | ((~c1)&(~c3)&(c4)&(~c6)) | ((c2)&(c3)&(c4)&(c6)) | ((c1)&(c3)&(c4)&(c6)) | ((c1)&(c2)&(c3)&(c6)) | ((c1)&(c2)&(c3)&(c4)) | ((c1)&(c2)&(c4)&(c6)));

assign D = (((~c1)&(~c2)&(~c3)&(~c4)&(~c6))| ((c1)&(c2)&(c3)&(c4)&(c6)) | ((c2)&(c3)&(~c4)&(~c6)) | ((~c1)&(~c2)&(c4)&(c6)) | ((~c1)&(c3)&(~c4)&(c6)) | ((~c1)&(c3)&(c4)&(~c6)) | ((c1)&(c2)&(~c3)&(~c4)) | ((c1)&(~c2)&(c3)&(~c4)) | ((c1)&(~c2)&(~c3)&(c6)) | ((c1)&(~c2)&(c4)&(~c6)) | ((c2)&(~c3)&(c4)&(~c6)));

assign E = (((~c1)&(c2)&(~c3)&(c4)&(c6)) | ((~c1)&(c2)&(c3)&(~c4)&(c6)) | ((~c1)&(~c2)&(c3)&(c4)&(c6)) | ((~c1)&(c2)&(c3)&(c4)&(~c6)) | ((c1)&(c2)&(c3)&(~c4)&(~c6)) | ((c1)&(c2)&(~c3)&(~c4)&(c6)) | ((c1)&(~c2)&(c3)&(~c4)&(c6)) | ((c1)&(~c2)&(~c3)&(c4)&(c6)) | ((c1)&(c2)&(c3)&(c4)&(c6)) | ((c1)&(~c2)&(c3)&(c4)&(~c6)) | ((c1)&(c2)&(~c3)&(c4)&(~c6)));

assign F = (((c1)&(c2)&(c3)&(c4)&(c6)) | ((~c2)&(~c3)&(~c4)&(~c6)) | ((~c1)&(~c2)&(~c3)&(~c4)) | ((~c1)&(~c2)&(~c4)&(~c6)) | ((~c1)&(~c2)&(~c3)&(c6)) | ((~c1)&(~c3)&(~c4)&(~c6)));

assign G = (((~c2)&(~c3)) | ((~c2)&(c3)&(~c4)) | ((~c1)&(c2)&(~c3)) | ((c2)&(~c3)&(~c4)) | ((c2)&(c3)&(~c4)&(~c6)) | ((~c1)&(c2)&(~c4)&(c6)) | ((~c1)&(~c2)&(c4)) | ((c2)&(~c3)&(c4)&(~c6)) | ((~c2)&(c4)&(~c6)) | ((~c1)&(c4)&(~c6)));

endmodule