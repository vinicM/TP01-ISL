module display (
    input C1,
    input C2,
    input C3,
    input C4,
    input C5,


    output A,
    output B,
    output C,
    output D
);
    
endmodule