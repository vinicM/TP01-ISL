module maquina (
    
    input 


);
    
endmodule