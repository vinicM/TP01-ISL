module display (

    input c1,
    input c2,
    input c3,
    input c4,
    input c5,

    output a,
    output b,
    output c,
    output d,
    output e,
    output f,
    output g
    
);

assign a = ((~c1) & (~c2) & c3 & c4)| ((~c1) & c2 & c4 & (~c5)) | ((~c2) & c3 & (~c4) & c5) | ((~c1) & c2 & (~c3) & c5) | (c1 & c3 & (~c4) & (~c5)) | (c1 & (~c2) & c4 & (~c5)) | (c1 & (~c3) &(~c4) & c5) | (c1 & c2 & (~c3) & (~c5)) | ((~c1) & c2 & c3 & (~c4)) | ((~c2) & (~c3) & c4 & c5) | (c1 & c2 & c3 & c4 & c5) | ((~c1) & (~c2) & (~c3) & (~c4) & (~c5));
assign b = (c5) | (c4) | (c3) | (c2) | (c1);
assign c = ((~c1) & (~c2) & (~c3)) | ((~c1) & (~c2) & (~c4)) | ((~c1) & (~c3) & (~c4)) | ((~c2) & (~c3) &(~c4)) | ((~c1) & (~c2) & (~c5)) | ((~c1) & (~c3) & (~c5)) | ((~c2) & (~c3) & (~c5)) | ((~c1) & (~c4) & (~c5)) | ((~c2) & (~c4) & (~c5)) | ((~c3) & (~c4) & (~c5)) | (c2 & c3 & c4 & c5) | (c1 & c3 & c4 & c5) | (c1 & c2 & c4 & c5) | (c1 & c2 & c3 & c5) | (c1 & c2 & c3 & c4);
assign d = ((~c1) & (~c2) & c4 & c5) | (c1 & c2 & (~c3) & (~c4)) | (c1 & (~c2) & (~c3) & c5) | ((~c1) & c3 & c4 & (~c5)) | (c2 & c3 & (~c4) & (~c5)) | ((~c1) & c3 & (~c4) & c5) | (c2 & (~c3) & c4 & (~c5)) | (c1 & (~c2) & c4 & (~c5)) | ((~c1) & c2 & (~c3) & c5) | (c1 & (~c2) & c3 & (~c4)) | (c1 & c2 & c3 & c4 & c5) | ((~c1) & (~c2) & (~c3) & (~c4) & (~c5));
assign e = ((~c1) & (~c2) & c3 & c4 & c5) | ((~c1) & c2 & (~c3) & c4 & c5) | ((~c1) & c2 & c3 & (~c4) & c5) | ((~c1) & c2 & c3 & c4 & (~c5)) | (c1 & (~c2) & (~c3) & c4 & c5) | (c1 & (~c2) & c3 & (~c4) & c5) | (c1 & (~c2) & c3 & c4 & (~c5)) | (c1 & c2 & (~c3) & (~c4) & c5) | (c1 & c2 & (~c3) & c4 & (~c5)) | (c1 & c2 & c3 & (~c4) & (~c5)) | (c1 & c2 & c3 & c4 & c5);
assign f = ((~c1) & (~c2) & (~c3) & (~c4)) | ((~c1) & (~c2) & (~c3) & (~c5)) | ((~c1) & (~c2) & (~c4) & (~c5)) | ((~c1) & (~c3) &(~c4) & (~c5)) | ((~c2) & (~c3) & (~c4) & (~c5)) | (c1 & c2 & c3 & c4 & c5);
assign g = ((~c1) & (~c2)) | ((~c1) & (~c3)) | ((~c2) & (~c3)) | ((~c1) & (~c4)) | ((~c2) & (~c4)) | ((~c3) & (~c4)) | ((~c1) & (~c5)) | ((~c2) & (~c5)) | ((~c3) & (~c5)) | ((~c4) & (~c5));


endmodule