module display (
    input c1,
    input c2,
    input c3,
    input c4,
    input c5,


    output A,
    output B,
    output C,
    output D,
    output E,
    output F,
    output G
);

assign A = (((~c1)&(c2)&(~c3)&(c5)) | ((~c1)&(c2)&(c3)&(~c4)) | ((~c1)&(c2)&(c4)&(~c5)) | ((~c1)&(~c2)&(c3)&(c4)) | ((~c1)&(~c2)&(~c3)&(~c4)&(~c5)) | ((~c1)&(~c2)&(~c3)&(~c4)&(c5)) | ((~c1)&(~c2)&(~c3)&(c4)&(c5)) | ((c1)&(c2)&(~c3)&(~c4)) | ((c1)&(c3)&(~c4)&(~c5)) | ((c1)&(~c2)&(c4)&(~c5)) | ((c1)&(~c2)&(~c3)&(c5)) | ((c1)&(c2)&(c3)&(c4)&(c5)) | ((c1)&(c2)&(~c3)&(c4)&(~c5)));
//assign A = (((~c1)&(~c2)&(~c3)&(~c4)&(~c5))| ((c1)&(c2)&(c3)&(c4)&(c5)) | ((c2)&(c3)&(~c4)&(~c5)) | ((~c1)&(~c2)&(c4)&(c5)) | ((~c1)&(c3)&(~c4)&(c5)) | ((~c1)&(c3)&(c4)&(~c5)) | ((c1)&(c2)&(~c3)&(~c4)) | ((c1)&(~c2)&(c3)&(~c4)) | ((c1)&(~c2)&(~c3)&(c5)) | ((c1)&(~c2)&(c4)&(~c5)) | ((c2)&(~c3)&(c4)&(~c5)) | ((c1)&(~c2)&(c4)&(~c5))));

assign B = ((c2) | ((~c2)&(c3)) | ((~c2)&(~c3)&(~c4)&(c5)) | ((~c2)&(~c3)&(c4)) | ((c1)&(~c2)&(~c3)&(~c4)&(~c5)));

assign C = (((~c2)&(~c4)&(~c5)) | ((~c1)&(~c4)&(~c5)) | ((~c2)&(~c3)&(~c4)&(c5)) | ((~c1)&(~c2)&(~c3)&(c5)) | ((~c1)&(~c2)&(c4)&(~c5)) | ((c1)&(~c2)&(~c3)&(~c4)) | ((c2)&(~c3)&(~c4)&(~c5)) | ((~c1)&(~c2)&(~c4)&(c5)) | ((~c1)&(~c3)&(~c4)&(c5)) | ((~c1)&(~c3)&(c4)&(~c5)) | ((c2)&(c3)&(c4)&(c5)) | ((c1)&(c3)&(c4)&(c5)) | ((c1)&(c2)&(c3)&(c5)) | ((c1)&(c2)&(c3)&(c4)) | ((c1)&(c2)&(c4)&(c5)));

assign D = (((~c1)&(c2)&(c3)&(~c4)&(~c5)) | ((~c1)&(c2)&(~c4)&(c5)) | ((~c1)&(c2)&(~c3)&( c4)) | ((~c1)&(c3)&(c4)&(~c5)) | ((~c1)&(~c2)&(c4)&(c5)) | ((~c1)&(~c2)&(c3)&(~c4)&(c5)) | ((~c1)&(~c2)&(~c3)&(~c4)&(~c5)) | ((c1)&(c2)&(~c3)&(~c4)) | ((c1)&(c3)&(~c4)&(c5)) | ((c1)&(~c2)&(~c4)&(c5)) | ((c1)&(~c2)&(~c3)&(c4)) | ((c1)&(~c2)&(c3)&(c4)&(~c5)) | ((c1)&(c2)&(c3)&(c4)&(c5)) | ((c1)&(c2)&(~c3)&(c4)&(~c5)));

//assign D = (((~c1)&(~c2)&(~c3)&(~c4)&(~c5))| ((c1)&(c2)&(c3)&(c4)&(c5)) | ((c2)&(c3)&(~c4)&(~c5)) | ((~c1)&(~c2)&(c4)&(c5)) | ((~c1)&(c3)&(~c4)&(c5)) | ((~c1)&(c3)&(c4)&(~c5)) | ((c1)&(c2)&(~c3)&(~c4)) | ((c1)&(~c2)&(c3)&(~c4)) | ((c1)&(~c2)&(~c3)&(c5)) | ((c1)&(~c2)&(c4)&(~c5)) | ((c2)&(~c3)&(c4)&(~c5)));

assign E = (((~c1)&(c2)&(~c3)&(c4)&(c5)) | ((~c1)&(c2)&(c3)&(~c4)&(c5)) | ((~c1)&(~c2)&(c3)&(c4)&(c5)) | ((~c1)&(c2)&(c3)&(c4)&(~c5)) | ((c1)&(c2)&(c3)&(~c4)&(~c5)) | ((c1)&(c2)&(~c3)&(~c4)&(c5)) | ((c1)&(~c2)&(c3)&(~c4)&(c5)) | ((c1)&(~c2)&(~c3)&(c4)&(c5)) | ((c1)&(c2)&(c3)&(c4)&(c5)) | ((c1)&(~c2)&(c3)&(c4)&(~c5)) | ((c1)&(c2)&(~c3)&(c4)&(~c5)));

assign F = (((~c1)&(c2)&(~c3)&(~c4)&(~c5)) | ((~c1)&(~c2)&(~c4)&(~c5)) | ((~c1)&(~c2)&(~c3)&(~c4)&(c5)) | ((~c1)&(~c2)&(~c3)&(c4)&(~c5)) | ((c1)&(c2)&(c3)&(c4)&(c5)) | ((c1)&(~c2)&(~c3)&(~c4)&(~c5)));
//assign F = (((c1)&(c2)&(c3)&(c4)&(c5)) | ((~c2)&(~c3)&(~c4)&(~c5)) | ((~c1)&(~c2)&(~c3)&(~c4)) | ((~c1)&(~c2)&(~c4)&(~c5)) | ((~c1)&(~c2)&(~c3)&(c5)) | ((~c1)&(~c3)&(~c4)&(~c5)));

assign G = (((~c2)&(~c3)) | ((~c2)&(c3)&(~c4)) | ((~c1)&(c2)&(~c3)) | ((c2)&(~c3)&(~c4)) | ((c2)&(c3)&(~c4)&(~c5)) | ((~c1)&(c2)&(~c4)&(c5)) | ((~c1)&(~c2)&(c4)) | ((c2)&(~c3)&(c4)&(~c5)) | ((~c2)&(c4)&(~c5)) | ((~c1)&(c4)&(~c5)));

endmodule