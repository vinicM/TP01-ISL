module ff(

    input data,
    input c,
    input r,
    output q;

);
endmodule

module maquina (
    
    input clk,
    input reset,
    output s1,
    output s2,


);
    
endmodule