module ff(

    input data,
    input c,
    input r,
    output q;

);
endmodule

module maquina (
    
    input clk,
    input reset,
    output saldoInsuf,
    output trocoRec,
    output doceComp,
    output doceEtroco;


);
    
endmodule